LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY Shameem_03132022_DFlipFlopMasterSlave IS 
	PORT (Shameem_03132022_D: IN STD_LOGIC;
		   Shameem_03132022_CLK: IN STD_LOGIC;
		   Shameem_03132022_PRN: IN STD_LOGIC;
		   Shameem_03132022_CLRN: IN STD_LOGIC;
		   Shameem_03132022_Q: OUT STD_LOGIC);
END Shameem_03132022_DFlipFlopMasterSlave;

ARCHITECTURE bdf_type OF Shameem_03132022_DFlipFlopMasterSlave IS 
SIGNAL  Shameem_03132022_SYNTHESIZED_WIRE_0,  Shameem_03132022_SYNTHESIZED_WIRE_1: STD_LOGIC;
BEGIN 
	PROCESS( Shameem_03132022_CLRN, Shameem_03132022_PRN, Shameem_03132022_SYNTHESIZED_WIRE_0, Shameem_03132022_D)
	BEGIN
		IF (Shameem_03132022_CLRN = '0') THEN
			Shameem_03132022_SYNTHESIZED_WIRE_1 <= '0';
		ELSIF (Shameem_03132022_PRN = '0') THEN
			Shameem_03132022_SYNTHESIZED_WIRE_1 <= '1';
		ELSIF (Shameem_03132022_SYNTHESIZED_WIRE_0 = '1') THEN
			Shameem_03132022_SYNTHESIZED_WIRE_1 <=  Shameem_03132022_D;
	END IF;
	END PROCESS;
	PROCESS( Shameem_03132022_CLRN, Shameem_03132022_PRN, Shameem_03132022_CLK, Shameem_03132022_SYNTHESIZED_WIRE_1)
	BEGIN
		IF (Shameem_03132022_CLRN = '0') THEN
			Shameem_03132022_Q <= '0';
		ELSIF (Shameem_03132022_PRN = '0') THEN
			Shameem_03132022_Q <= '1';
		ELSIF (Shameem_03132022_CLK = '1') THEN
			Shameem_03132022_Q <= Shameem_03132022_SYNTHESIZED_WIRE_1;
	END IF;
	END PROCESS;
Shameem_03132022_SYNTHESIZED_WIRE_0 <= NOT(Shameem_03132022_CLK);
END bdf_type;